`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author:Niculescu Vlad
// Module Name:    Transcoder 
//////////////////////////////////////////////////////////////////////////////////
module Transcoder ( output reg[15:0] out,
input [3:0] in
);

always@(*) begin
case(in)
4'd0: out[15:0] = 16'b0000000000000000;
4'd1: out[15:0] = 16'b0000000000000010;
4'd2: out[15:0] = 16'b0000000000000100;
4'd3: out[15:0] = 16'b0000000000001000;
4'd4: out[15:0] = 16'b0000000000010000;
4'd5: out[15:0] = 16'b0000000000100000;
4'd6: out[15:0] = 16'b0000000001000000;
4'd7: out[15:0] = 16'b0000000010000000;
4'd8: out[15:0] = 16'b0000000100000000;
4'd9: out[15:0] = 16'b0000001000000000;
4'hA: out[15:0] = 16'b0000010000000000;
4'hB: out[15:0] = 16'b0000100000000000;
4'hC: out[15:0] = 16'b0001000000000000;
4'hD: out[15:0] = 16'b0010000000000000;
4'hE: out[15:0] = 16'b0100000000000000;
4'hF: out[15:0] = 16'b1111111111111111;
endcase
end
endmodule