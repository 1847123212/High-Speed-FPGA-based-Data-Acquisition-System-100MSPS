`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
// Author:Niculescu Vlad
// Module Name:    Square 
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module Square(a,b,p
    );
input  [9:0]  a;
input  [9:0]  b;
output [19:0] p;
mult your_instance_name (
  .a(a), // input [9 : 0] a
  .b(b), // input [9 : 0] b
  .p(p) // output [19 : 0] p
);
endmodule
