`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Author:Niculescu Vlad
// Module Name:    MUX 
//////////////////////////////////////////////////////////////////////////////////
module MUX(input [10:0] a, input [10:0] b, input sel, output [10:0] out
    );

assign out = sel ? a : b;
endmodule
