`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author:Niculescu Vlad
// Module Name:    MUX_converter 
//////////////////////////////////////////////////////////////////////////////////
module MUX_converter(input [8:0] a, input sel, output [8:0] x
    );

assign x = sel ? a : ~a + 1;

endmodule
