--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package defs is

type slv8array is array (natural range <>) of std_logic_vector(7 downto 0);

end defs;

package body defs is

end defs;
